module Part3(input logic [2:0]in, output logic [1:0]out);
	FullAdder FA(in);
endmodule