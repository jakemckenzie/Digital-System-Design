module Mux_3w_5_to_1(input S0,S1,S2,input [2:0]u,v,w,x,y,output [2:0]m);
   assign w0 = S0 ? v : u;
   assign w1 = S0 ? x : w;
   assign w2 = S1 ? w1 : w0;
   assign m = S2 ? y : w2;
endmodule // Mux_3w_5_to_1

module Mux_3w_5_to_1_testbench();
   reg [2:0]u,v,w,x,y;
   reg S0,S1,S2;
   wire [2:0] m;

   Mux_3w_5_to_1 DUT(S0,S1,S2,u,v,w,x,y,m);
   initial begin
		u = 1; v = 2;w = 3;x = 4;y = 5;
      S0 = 0;S1 = 0;S2 = 0;#10;
      S0 = 1;S1 = 0;S2 = 0;#10;
      S0 = 0;S1 = 1;S2 = 0;#10;
      S0 = 1;S1 = 1;S2 = 0;#10;
      S0 = 0;S1 = 0;S2 = 1;#10;
   end

endmodule // Mux_3w_5_to_1_testbench
