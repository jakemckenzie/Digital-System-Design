Epimetheus@EPIMETHEUS-PC.18312:1522626642