module Part2();

endmodule