module notes_4_18();
    //read the book, the examples weren't reproducible because she started with existing code
endmodule