module Part5([17:0]SW);
    input [17:0]SW;
    output [0:6]Hex;

    always @(*)
    begin
        case(C)
        always @(*)
            begin
                case(SW[14:12])
            end
        always @(*)
            begin
                case(SW[11:9)
            end
        always @(*)
            begin
                case(SW[8:6)
            end
        always @(*)
            begin
                case(SW[5:3)
            end
    end
endmodule

//ask about big endian vs little endian for input vs output
//use more asserts
//always put a $stop

//display = print
//monitor is printf

//You typically do things little endian