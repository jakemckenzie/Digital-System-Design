module Decode_part2();

endmodule