//TCES330 Spring 2018
//Using LPMs examples
//This module includes an Altera LPM adder
//J. Sheng

module TestLPM3(A,B,Cin,S,Cout);

	input [15:0]A,B;
	input Cin;
	output [15:0]S;
	output Cout;

	AlteraAdder MyAdder1(
	.cin(Cin),
	.dataa(A),
	.datab(B),
	.cout(Cout),
	.result(S));

endmodule


///
`timescale 1ps/1ps
module TestLPM3_testbench();

	logic [15:0]A,B;
	logic Cin;
	logic [15:0]S;
	logic Cout;

	TestLPM3 DUT (A,B,Cin,S,Cout);

	integer I;

	initial begin
		Cin=0;
		for (I=0; I<50; I++) begin
			A=$urandom;
			B=$urandom;
			Cin=1;
			assert ({Cout,S} == A+B+Cin);

			#10;
			Cin=0;
			assert ({Cout,S} == A+B+Cin);
			#10;
			A=$urandom;
			B=$urandom;
			Cin=0;
			assert ({Cout,S} == A+B+Cin);

			#10;
			Cin=1;
			assert ({Cout,S} == A+B+Cin);
			#10;
		end
	$stop;
	end
	
	initial begin
		$monitor ($time,,,A,,,B,,,Cin,,,{Cout, S});
	end


endmodule
