module notes_4_18();

endmodule